module regfile( 
    ctrl_bus_if.central ctrl_bus,
    input   logic[5:0]  reg_num,
);
    
endmodule
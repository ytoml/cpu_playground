module hazard_unit(
	input	logic		rs_E, rt_E, rd_E,
	input	logic[4:0]	reg_id_M, reg_id_W,
	input	logic		reg_write_M, reg_write_W,
	output	logic		forwardA_E, forwardB_E
);
	// TODO
endmodule
`include "lib_cpu.svh"
module decoder import lib_cpu::*;(
    mem_bus_if.central  imem_bus,
    output  OPECODE     op,
    output  FUNCT       funct
);

    
endmodule
module datapath(
    ctrl_bus_if.central ctrl_bus
);
    sign_ext    sign_ext();
    alu         alu();
    
endmodule
module datapath(
    ctrl_bus_if.central ctrl_bus
);
    
endmodule